`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2019/05/15 18:23:15
// Design Name:
// Module Name: vga_param
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

/* VGA(640?��~480)?��p?��?��?��?��?��[?��^ */
localparam WHITE   = 3'b000;
localparam BLACK   = 3'b001;
localparam RED     = 3'b010;
localparam BLUE    = 3'b011;
localparam GREEN   = 3'b100;
localparam YELLOW  = 3'b101;
localparam LIGHTB  = 3'b110;
localparam PINK    = 3'b111;