`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/05/27 18:35:20
// Design Name: 
// Module Name: adau1761_configuraiton_data
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adau1761_configuraiton_data(
    input               clk,
    input      [9:0]    address,
    output reg [8:0]    data
    );
    
    always @(posedge clk) begin
        case(address)
        10'b0000000000: data <= 9'b011101111;
        10'b0000000001: data <= 9'b101110110;//1:I2S START R0���W�X�^�iClock control�j��1110����� INFREQ[1:0] = 1024*fs core clock desenable
        10'b0000000010: data <= 9'b101000000;
        10'b0000000011: data <= 9'b100000000;
        10'b0000000100: data <= 9'b100001110;
        10'b0000000101: data <= 9'b011111111; //I2S STOP
        10'b0000000110: data <= 9'b101110110; //2:I2S START R1���W�X�^�iPLL control�j�� 
        10'b0000000111: data <= 9'b101000000;
        10'b0000001000: data <= 9'b100000010;
        10'b0000001001: data <= 9'b100000000; //�����ȍ~�̐��l���Ԃ�����
        10'b0000001010: data <= 9'b101111101; //00000000,01111101,00000000,00001100,00100011,00000001 M=125 X=2 R=4 N=12 Mode=512*48k = 24.576MHz
        10'b0000001011: data <= 9'b100000000; //48kHz�œ���!
        10'b0000001100: data <= 9'b100001100;
        10'b0000001101: data <= 9'b100100011; //X:01 = X=2
        10'b0000001110: data <= 9'b100000001;//PLL enable
        10'b0000001111: data <= 9'b011111111;//I2S STOP
        10'b0000010000: data <= 9'b011101111;//delay PLL rock���Ԋm��
        10'b0000010001: data <= 9'b101110110;//3:I2S START R0���W�X�^�iClock control�j��1111����� core clock enable
        10'b0000010010: data <= 9'b101000000;
        10'b0000010011: data <= 9'b100000000;
        10'b0000010100: data <= 9'b100001111;
        10'b0000010101: data <= 9'b011111111;//4:I2S STOP
        10'b0000010110: data <= 9'b011101111;//delay
        10'b0000010111: data <= 9'b101110110;//5:I2S START R15�iSerial Port 0�j��1����� ���g��fs��I2c mode �ŃN���b�N���}�X�^�[�ɑ����Ă����
        10'b0000011000: data <= 9'b101000000;
        10'b0000011001: data <= 9'b100010101;
        10'b0000011010: data <= 9'b100000001;
        10'b0000011011: data <= 9'b011111111;//I2S STOP
        10'b0000011100: data <= 9'b101110110;//6:I2S START R10�iRecord mic bias�j��1����� ebable
        10'b0000011101: data <= 9'b101000000;
        10'b0000011110: data <= 9'b100001010;
        10'b0000011111: data <= 9'b100000001;
        10'b0000100000: data <= 9'b011111111;//I2S STOP
        10'b0000100001: data <= 9'b101110110;//7:I2S START R11�iALC 0�j��5����� ALC�͉��̐ݒ�ɕK�v
        10'b0000100010: data <= 9'b101000000;
        10'b0000100011: data <= 9'b100001011;
        10'b0000100100: data <= 9'b100000101;
        10'b0000100101: data <= 9'b011111111;//I2S STOP
        10'b0000100110: data <= 9'b101110110;//8:I2S START R12�iALC 1�j��1�����
        10'b0000100111: data <= 9'b101000000;
        10'b0000101000: data <= 9'b100001100;
        10'b0000101001: data <= 9'b100000001;
        10'b0000101010: data <= 9'b011111111;//I2S STOP
        10'b0000101011: data <= 9'b101110110;//9:I2S START R13�iALC 2�j��5�����
        10'b0000101100: data <= 9'b101000000;
        10'b0000101101: data <= 9'b100001101;
        10'b0000101110: data <= 9'b100000101;
        10'b0000101111: data <= 9'b011111111;//I2S STOP
        10'b0000110000: data <= 9'b101110110;//10:I2S START R22�iPlay Mixer Left 0�j33�����
        10'b0000110001: data <= 9'b101000000;
        10'b0000110010: data <= 9'b100011100;
        10'b0000110011: data <= 9'b100100001;
        10'b0000110100: data <= 9'b011111111;//I2S STOP
        10'b0000110101: data <= 9'b101110110;//11:I2S START R24�iPlay Mixer Right 0�j��65�����
        10'b0000110110: data <= 9'b101000000;
        10'b0000110111: data <= 9'b100011110;
        10'b0000111000: data <= 9'b101000001;
        10'b0000111001: data <= 9'b011111111;//I2S STOP
        10'b0000111010: data <= 9'b101110110;//12:I2S START  R29�iPlay HP left vol�j��231����
        10'b0000111011: data <= 9'b101000000;
        10'b0000111100: data <= 9'b100100011;
        10'b0000111101: data <= 9'b111100111;
        10'b0000111110: data <= 9'b011111111;//I2S STOP
        10'b0000111111: data <= 9'b101110110;//13:I2S START R30�iPlay HP right vol�j��231����
        10'b0001000000: data <= 9'b101000000;
        10'b0001000001: data <= 9'b100100100;
        10'b0001000010: data <= 9'b111100111;
        10'b0001000011: data <= 9'b011111111;//I2S STOP
        10'b0001000100: data <= 9'b101110110;//14:I2S START R31�iLine output left vol�j��231����
        10'b0001000101: data <= 9'b101000000;
        10'b0001000110: data <= 9'b100100101;
        10'b0001000111: data <= 9'b111100111;
        10'b0001001000: data <= 9'b011111111;//I2S STOP
        10'b0001001001: data <= 9'b101110110;//15:I2S START R32�iLine output right vol�j��231����
        10'b0001001010: data <= 9'b101000000;
        10'b0001001011: data <= 9'b100100110;
        10'b0001001100: data <= 9'b111100111;
        10'b0001001101: data <= 9'b011111111;//I2S STOP
        10'b0001001110: data <= 9'b101110110;//16:I2S START R19�iADC control�j��3����
        10'b0001001111: data <= 9'b101000000;
        10'b0001010000: data <= 9'b100011001;
        10'b0001010001: data <= 9'b100000011;
        10'b0001010010: data <= 9'b011111111;//I2S STOP
        10'b0001010011: data <= 9'b101110110;//17:I2S START R35�iPlay power mgmt�j��3����
        10'b0001010100: data <= 9'b101000000;
        10'b0001010101: data <= 9'b100101001;
        10'b0001010110: data <= 9'b100000011;
        10'b0001010111: data <= 9'b011111111;//I2S STOP
        10'b0001011000: data <= 9'b101110110;//18:I2S START R36�iDAC Control 0�j��3����
        10'b0001011001: data <= 9'b101000000;
        10'b0001011010: data <= 9'b100101010;
        10'b0001011011: data <= 9'b100000011;
        10'b0001011100: data <= 9'b011111111;//I2S STOP
        10'b0001011101: data <= 9'b101110110;//19:I2S START R58�iSerial input routecontrol�j��1����
        10'b0001011110: data <= 9'b101000000;
        10'b0001011111: data <= 9'b111110010;
        10'b0001100000: data <= 9'b100000001;
        10'b0001100001: data <= 9'b011111111;//I2S STOP
        10'b0001100010: data <= 9'b101110110;//20:I2S START R59�iSerial output routecontrol�j��1����
        10'b0001100011: data <= 9'b101000000;
        10'b0001100100: data <= 9'b111110011;
        10'b0001100101: data <= 9'b100000001;
        10'b0001100110: data <= 9'b011111111;//I2S STOP
        10'b0001100111: data <= 9'b101110110;//21:I2S START R65�iClock Enable 0�j��127����
        10'b0001101000: data <= 9'b101000000;
        10'b0001101001: data <= 9'b111111001;
        10'b0001101010: data <= 9'b101111111;
        10'b0001101011: data <= 9'b011111111;//I2S STOP
        10'b0001101100: data <= 9'b101110110;//22:I2S START R66�iClock Enable 1�j��3����
        10'b0001101101: data <= 9'b101000000;
        10'b0001101110: data <= 9'b111111010;
        10'b0001101111: data <= 9'b100000011;
        10'b0001110000: data <= 9'b011111111;//I2S STOP
        10'b0001110001: data <= 9'b000010011;//JUMP pc <= 0010011000 pc = 114
        10'b0010011000: data <= 9'b010000000;//�ݒ肪�I������炱���ɗ��� skip_clear skip = 1 pc = 152
        10'b0010011001: data <= 9'b000010100;//JUMP pc <= 0010100000 skip
        10'b0010011010: data <= 9'b010000001;//skip clear skip = 1
        10'b0010011011: data <= 9'b000011001;//JUMP pc <= 0011001000 skip
        10'b0010011100: data <= 9'b000010011;//JUMP pc <= 0010011000
        default       : data <= 9'b010000000; 
        endcase
    end
    
endmodule
