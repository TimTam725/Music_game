`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/06/01 00:34:21
// Design Name: 
// Module Name: audio_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module audio_mem(
//    input                clk,
//    input                rst,
    input      [8:0]     pc,
    output     [8:0]     data
    );
    
    assign data = (pc == 9'd0)  ?  {5'd0,  4'd15} ://0�@
                   (pc == 9'd1)  ?  {5'd17, 4'd1} :
                   (pc == 9'd2)  ?  {5'd17, 4'd1} :
                   (pc == 9'd3)  ?  {5'd0,  4'd1} :
                   (pc == 9'd4)  ?  {5'd17, 4'd1} :
                   (pc == 9'd5)  ?  {5'd0 , 4'd1} :
                   (pc == 9'd6)  ?  {5'd13, 4'd1} :
                   (pc == 9'd7)  ?  {5'd17, 4'd1} :
                   (pc == 9'd8)  ?  {5'd0,  4'd1} ://1�@�~�~�E�~�E�h�~�E
                   (pc == 9'd9)  ?  {5'd20, 4'd1} :
                   (pc == 9'd10) ?  {5'd0,  4'd5} :
                   (pc == 9'd11) ?  {5'd8,  4'd1} :
                   (pc == 9'd12) ?  {5'd0,  4'd5} ://2�@�\�E�E�E�\�E�E�E
                   (pc == 9'd13) ?  {5'd13,  4'd1} :
                   (pc == 9'd14) ?  {5'd0,  4'd3} :
                   (pc == 9'd15) ?  {5'd8,  4'd1} :
                   (pc == 9'd16) ?  {5'd0,  4'd3} :
                   (pc == 9'd17) ?  {5'd5,  4'd1} ://3�@�h�E�E�E�\�E�E�E�~
                   (pc == 9'd18) ?  {5'd0,  4'd3} :
                   (pc == 9'd19) ?  {5'd10,  4'd1} :
                   (pc == 9'd20) ?  {5'd0,  4'd1} :
                   (pc == 9'd21) ?  {5'd12,  4'd1} :
                   (pc == 9'd22) ?  {5'd0,  4'd1} :
                   (pc == 9'd23) ?  {5'd11,  4'd1} :
                   (pc == 9'd24) ?  {5'd10,  4'd1} :
                   (pc == 9'd25) ?  {5'd0,  4'd1} ://4�@�E�E�E���E�V�E�V���E
                   (pc == 9'd26) ?  {5'd8,  4'd2} :
                   (pc == 9'd27) ?  {5'd17,  4'd2} :
                   (pc == 9'd28) ?  {5'd20,  4'd1} :
                   (pc == 9'd29) ?  {5'd23,  4'd1} :
                   (pc == 9'd30) ?  {5'd0,  4'd1} :
                   (pc == 9'd31) ?  {5'd18,  4'd1} :
                   (pc == 9'd32) ?  {5'd20,  4'd1} : //5�@�\�~�\���E�t�@�\
                   (pc == 9'd33) ?  {5'd0,  4'd1} :
                   (pc == 9'd34) ?  {5'd17,  4'd1} :
                   (pc == 9'd35) ?  {5'd0,  4'd1} :
                   (pc == 9'd36) ?  {5'd13,  4'd1} :
                   (pc == 9'd37) ?  {5'd15,  4'd1} :
                   (pc == 9'd38) ?  {5'd12,  4'd1} :
                   (pc == 9'd39) ?  {5'd0,  4'd3} : //6�@�E�~�E�h���V�E�E�E
                   (pc == 9'd40) ?  {5'd13,  4'd1} :
                   (pc == 9'd41) ?  {5'd0,  4'd3} :
                   (pc == 9'd42) ?  {5'd8,  4'd1} :
                   (pc == 9'd43) ?  {5'd0,  4'd3} :
                   (pc == 9'd44) ?  {5'd5,  4'd1} ://7�@�h�E�E�E�\�E�E�E�~ (�Q�T��)
                   (pc == 9'd45) ?  {5'd0,  4'd3} :
                   (pc == 9'd46) ?  {5'd10,  4'd1} :
                   (pc == 9'd47) ?  {5'd0,  4'd1} :
                   (pc == 9'd48) ?  {5'd12,  4'd1} :
                   (pc == 9'd49) ?  {5'd0,  4'd1} :
                   (pc == 9'd50) ?  {5'd11,  4'd1} :
                   (pc == 9'd51) ?  {5'd10,  4'd1} :
                   (pc == 9'd52) ?  {5'd0,  4'd1} ://8�@�E�E�E���E�V�E�V���E
                   (pc == 9'd53) ?  {5'd8,  4'd2} :
                   (pc == 9'd54) ?  {5'd17,  4'd2} :
                   (pc == 9'd55) ?  {5'd20,  4'd1} :
                   (pc == 9'd56) ?  {5'd23,  4'd1} :
                   (pc == 9'd57) ?  {5'd0,  4'd1} :
                   (pc == 9'd58) ?  {5'd18,  4'd1} :
                   (pc == 9'd59) ?  {5'd20,  4'd1} ://9�@�\�~�\���E�t�@�\
                   (pc == 9'd60) ?  {5'd0,  4'd1} :
                   (pc == 9'd61) ?  {5'd17,  4'd1} :
                   (pc == 9'd62) ?  {5'd0,  4'd1} :
                   (pc == 9'd63) ?  {5'd13,  4'd1} :
                   (pc == 9'd64) ?  {5'd15,  4'd1} :
                   (pc == 9'd65) ?  {5'd12,  4'd1} :
                   (pc == 9'd66) ?  {5'd0,  4'd3} : //10�@�E�~�E�h���V�E�E�E (�Q�T�ڏI��)
                   (pc == 9'd67) ?  {5'd0,  4'd3} :
                   (pc == 9'd68) ?  {5'd20,  4'd1} :
                   (pc == 9'd69) ?  {5'd19,  4'd1} :
                   (pc == 9'd70) ?  {5'd18,  4'd1} :
                   (pc == 9'd71) ?  {5'd16,  4'd1} :
                   (pc == 9'd72) ?  {5'd0,  4'd1} :
                   (pc == 9'd73) ?  {5'd17,  4'd1} ://11�@�E�E�E�\�t�@�t�@���E�~
                   (pc == 9'd74) ?  {5'd0,  4'd1} :
                   (pc == 9'd75) ?  {5'd9,  4'd1} :
                   (pc == 9'd76) ?  {5'd10,  4'd1} :
                   (pc == 9'd77) ?  {5'd13,  4'd1} :
                   (pc == 9'd78) ?  {5'd0,  4'd1} :
                   (pc == 9'd79) ?  {5'd10,  4'd1} :
                   (pc == 9'd80) ?  {5'd13,  4'd1} :
                   (pc == 9'd81) ?  {5'd15,  4'd1} ://12�@�E�\���h�D���h��
                   (pc == 9'd82) ?  {5'd0,  4'd3} :
                   (pc == 9'd83) ?  {5'd20,  4'd1} :
                   (pc == 9'd84) ?  {5'd19,  4'd1} :
                   (pc == 9'd85) ?  {5'd18,  4'd1} :
                   (pc == 9'd86) ?  {5'd16,  4'd1} :
                   (pc == 9'd87) ?  {5'd0,  4'd1} :
                   (pc == 9'd88) ?  {5'd17,  4'd1} ://13�@�E�E�E�\�t�@�t�@���E�~
                   (pc == 9'd89) ?  {5'd0,  4'd1} :
                   (pc == 9'd90) ?  {5'd26,  4'd1} :
                   (pc == 9'd91) ?  {5'd0,  4'd1} :
                   (pc == 9'd92) ?  {5'd26,  4'd1} :
                   (pc == 9'd93) ?  {5'd26,  4'd1} :
                   (pc == 9'd94) ?  {5'd0,  4'd5} ://14�@�E�h�E�h�h�E�E�E�E�E�E
                   (pc == 9'd95) ?  {5'd0,  4'd3} :
                   (pc == 9'd96) ?  {5'd20,  4'd1} :
                   (pc == 9'd97) ?  {5'd19,  4'd1} :
                   (pc == 9'd98) ?  {5'd18,  4'd1} :
                   (pc == 9'd99) ?  {5'd16,  4'd1} :
                   (pc == 9'd100) ?  {5'd0,  4'd1} :
                   (pc == 9'd101) ?  {5'd17,  4'd1} ://15�@�E�E�E�\�t�@�t�@���E�~
                   (pc == 9'd102) ?  {5'd0,  4'd1} :
                   (pc == 9'd103) ?  {5'd9,  4'd1} :
                   (pc == 9'd104) ?  {5'd10,  4'd1} :
                   (pc == 9'd105) ?  {5'd13,  4'd1} :
                   (pc == 9'd106) ?  {5'd0,  4'd1} :
                   (pc == 9'd107) ?  {5'd10,  4'd1} :
                   (pc == 9'd108) ?  {5'd13,  4'd1} :
                   (pc == 9'd109) ?  {5'd15,  4'd1} ://16�@�E�\���h�D���h��
                   (pc == 9'd110) ?  {5'd0,  4'd3} :
                   (pc == 9'd111) ?  {5'd16,  4'd1} :
                   (pc == 9'd112) ?  {5'd0,  4'd3} :
                   (pc == 9'd113) ?  {5'd15,  4'd1} :
                   (pc == 9'd114) ?  {5'd0,  4'd3} ://17�@�~��
                   (pc == 9'd115) ?  {5'd13,  4'd1} :
                   (pc == 9'd116) ?  {5'd0,  4'd13} ://18�@�h�E�E�E
                   (pc == 9'd117) ?  {5'd0,  4'd3} :
                   (pc == 9'd118) ?  {5'd20,  4'd1} :
                   (pc == 9'd119) ?  {5'd19,  4'd1} :
                   (pc == 9'd120) ?  {5'd18,  4'd1} :
                   (pc == 9'd121) ?  {5'd16,  4'd1} :
                   (pc == 9'd122) ?  {5'd0,  4'd1} :
                   (pc == 9'd123) ?  {5'd17,  4'd1} ://19�@�E�E�E�\�t�@�t�@���E�~ (2�T��)
                   (pc == 9'd124) ?  {5'd0,  4'd1} :
                   (pc == 9'd125) ?  {5'd9,  4'd1} :
                   (pc == 9'd126) ?  {5'd10,  4'd1} :
                   (pc == 9'd127) ?  {5'd13,  4'd1} :
                   (pc == 9'd128) ?  {5'd0,  4'd1} :
                   (pc == 9'd129) ?  {5'd10,  4'd1} :
                   (pc == 9'd130) ?  {5'd13,  4'd1} :
                   (pc == 9'd131) ?  {5'd15,  4'd1} ://20�@�E�\���h�D���h��
                   (pc == 9'd132) ?  {5'd0,  4'd3} :
                   (pc == 9'd133) ?  {5'd20,  4'd1} :
                   (pc == 9'd134) ?  {5'd19,  4'd1} :
                   (pc == 9'd135) ?  {5'd18,  4'd1} :
                   (pc == 9'd136) ?  {5'd16,  4'd1} :
                   (pc == 9'd137) ?  {5'd0,  4'd1} :
                   (pc == 9'd138) ?  {5'd17,  4'd1} ://21�@�E�E�E�\�t�@�t�@���E�~
                   (pc == 9'd139) ?  {5'd0,  4'd1} :
                   (pc == 9'd140) ?  {5'd26,  4'd1} :
                   (pc == 9'd141) ?  {5'd0,  4'd1} :
                   (pc == 9'd142) ?  {5'd26,  4'd1} :
                   (pc == 9'd143) ?  {5'd26,  4'd1} :
                   (pc == 9'd144) ?  {5'd0,  4'd5} ://22�@�E�h�E�h�h�E�E�E�E�E�E
                   (pc == 9'd145) ?  {5'd0,  4'd3} :
                   (pc == 9'd146) ?  {5'd20,  4'd1} :
                   (pc == 9'd147) ?  {5'd19,  4'd1} :
                   (pc == 9'd148) ?  {5'd18,  4'd1} :
                   (pc == 9'd149) ?  {5'd16,  4'd1} :
                   (pc == 9'd150) ?  {5'd0,  4'd1} :
                   (pc == 9'd151) ?  {5'd17,  4'd1} ://23�@�E�E�E�\�t�@�t�@���E�~
                   (pc == 9'd152) ?  {5'd0,  4'd1} :
                   (pc == 9'd153) ?  {5'd9,  4'd1} :
                   (pc == 9'd154) ?  {5'd10,  4'd1} :
                   (pc == 9'd155) ?  {5'd13,  4'd1} :
                   (pc == 9'd156) ?  {5'd0,  4'd1} :
                   (pc == 9'd157) ?  {5'd10,  4'd1} :
                   (pc == 9'd158) ?  {5'd13,  4'd1} :
                   (pc == 9'd159) ?  {5'd15,  4'd1} ://24�@�E�\���h�D���h��
                   (pc == 9'd160) ?  {5'd0,  4'd3} :
                   (pc == 9'd161) ?  {5'd16,  4'd1} :
                   (pc == 9'd162) ?  {5'd0,  4'd3} :
                   (pc == 9'd163) ?  {5'd15,  4'd1} :
                   (pc == 9'd164) ?  {5'd0,  4'd3} ://25�@�~��
                   (pc == 9'd165) ?  {5'd13,  4'd1} :
                   (pc == 9'd166) ?  {5'd0,  4'd13} : //26�@�h
                   (pc == 9'd167) ?  {5'd13,  4'd1} :
                   (pc == 9'd168) ?  {5'd13,  4'd1} :
                   (pc == 9'd169) ?  {5'd0,  4'd1} :
                   (pc == 9'd170) ?  {5'd13,  4'd1} :
                   (pc == 9'd171) ?  {5'd0,  4'd1} :
                   (pc == 9'd172) ?  {5'd13,  4'd1} :
                   (pc == 9'd173) ?  {5'd15,  4'd1} :
                   (pc == 9'd174) ?  {5'd0,  4'd1} ://27�@�h�h�E�h�E�h��
                   (pc == 9'd175) ?  {5'd17,  4'd1} :
                   (pc == 9'd176) ?  {5'd13,  4'd1} :
                   (pc == 9'd177) ?  {5'd0,  4'd1} :
                   (pc == 9'd178) ?  {5'd10,  4'd1} :
                   (pc == 9'd179) ?  {5'd8,  4'd1} :
                   (pc == 9'd180) ?  {5'd0,  4'd5} ://28�@�~�h���\
                   (pc == 9'd181) ?  {5'd13,  4'd1} :
                   (pc == 9'd182) ?  {5'd13,  4'd1} :
                   (pc == 9'd183) ?  {5'd0,  4'd1} :
                   (pc == 9'd184) ?  {5'd13,  4'd1} :
                   (pc == 9'd185) ?  {5'd0,  4'd1} :
                   (pc == 9'd186) ?  {5'd13,  4'd1} :
                   (pc == 9'd187) ?  {5'd15,  4'd1} :
                   (pc == 9'd188) ?  {5'd17,  4'd1} ://29�@�h�h�E�h�E�h���~
                   (pc == 9'd189) ?  {5'd0,  4'd15} ://30�@�E�E�E
                   (pc == 9'd190) ?  {5'd13,  4'd1} :
                   (pc == 9'd191) ?  {5'd13,  4'd1} :
                   (pc == 9'd192) ?  {5'd0,  4'd1} :
                   (pc == 9'd193) ?  {5'd13,  4'd1} :
                   (pc == 9'd194) ?  {5'd0,  4'd1} :
                   (pc == 9'd195) ?  {5'd13,  4'd1} :
                   (pc == 9'd196) ?  {5'd15,  4'd1} :
                   (pc == 9'd197) ?  {5'd0,  4'd1} ://31�@�h�h�E�h�E�h��
                   (pc == 9'd198) ?  {5'd17,  4'd1} :
                   (pc == 9'd199) ?  {5'd13,  4'd1} :
                   (pc == 9'd200) ?  {5'd0,  4'd1} :
                   (pc == 9'd201) ?  {5'd10,  4'd1} :
                   (pc == 9'd202) ?  {5'd8,  4'd1} :
                   (pc == 9'd203) ?  {5'd0,  4'd5} ://32�@�~�h���\
                   (pc == 9'd204)  ?  {5'd17, 4'd1} :
                   (pc == 9'd205)  ?  {5'd17, 4'd1} :
                   (pc == 9'd206)  ?  {5'd0,  4'd1} :
                   (pc == 9'd207)  ?  {5'd17, 4'd1} :
                   (pc == 9'd208)  ?  {5'd0 , 4'd1} :
                   (pc == 9'd209)  ?  {5'd13, 4'd1} :
                   (pc == 9'd210)  ?  {5'd17, 4'd1} :
                   (pc == 9'd211)  ?  {5'd0,  4'd1} ://33�@�~�~�E�~�E�h�~�E
                   (pc == 9'd212)  ?  {5'd20, 4'd1} :
                   (pc == 9'd213) ?  {5'd0,  4'd5} :
                   (pc == 9'd214) ?  {5'd8,  4'd1} :
                   (pc == 9'd215) ?  {5'd0,  4'd5} ://34�@�\�E�E�E�\�E�E�E
                   (pc == 9'd216) ?  {5'd13,  4'd1} :
                   (pc == 9'd217) ?  {5'd0,  4'd3} :
                   (pc == 9'd218) ?  {5'd8,  4'd1} :
                   (pc == 9'd219) ?  {5'd0,  4'd3} :
                   (pc == 9'd220) ?  {5'd5,  4'd1} ://35�@�h�E�E�E�\�E�E�E�~
                   (pc == 9'd221) ?  {5'd0,  4'd3} :
                   (pc == 9'd222) ?  {5'd10,  4'd1} :
                   (pc == 9'd223) ?  {5'd0,  4'd1} :
                   (pc == 9'd224) ?  {5'd12,  4'd1} :
                   (pc == 9'd225) ?  {5'd0,  4'd1} :
                   (pc == 9'd226) ?  {5'd11,  4'd1} :
                   (pc == 9'd227) ?  {5'd10,  4'd1} :
                   (pc == 9'd228) ?  {5'd0,  4'd1} ://36�@�E�E�E���E�V�E�V���E
                   (pc == 9'd229) ?  {5'd8,  4'd2} :
                   (pc == 9'd230) ?  {5'd17,  4'd2} :
                   (pc == 9'd231) ?  {5'd20,  4'd1} :
                   (pc == 9'd232) ?  {5'd23,  4'd1} :
                   (pc == 9'd233) ?  {5'd0,  4'd1} :
                   (pc == 9'd234) ?  {5'd18,  4'd1} :
                   (pc == 9'd235) ?  {5'd20,  4'd1} : //37�@�\�~�\���E�t�@�\
                   (pc == 9'd236) ?  {5'd0,  4'd1} :
                   (pc == 9'd237) ?  {5'd17,  4'd1} :
                   (pc == 9'd238) ?  {5'd0,  4'd1} :
                   (pc == 9'd239) ?  {5'd13,  4'd1} :
                   (pc == 9'd240) ?  {5'd15,  4'd1} :
                   (pc == 9'd241) ?  {5'd12,  4'd1} :
                   (pc == 9'd242) ?  {5'd0,  4'd3} : //38�@�E�~�E�h���V�E�E�E
                   (pc == 9'd243) ?  {5'd13,  4'd1} :
                   (pc == 9'd244) ?  {5'd0,  4'd3} :
                   (pc == 9'd245) ?  {5'd8,  4'd1} :
                   (pc == 9'd246) ?  {5'd0,  4'd3} :
                   (pc == 9'd247) ?  {5'd5,  4'd1} ://39�@�h�E�E�E�\�E�E�E�~ (�Q�T��)
                   (pc == 9'd248) ?  {5'd0,  4'd3} :
                   (pc == 9'd249) ?  {5'd10,  4'd1} :
                   (pc == 9'd250) ?  {5'd0,  4'd1} :
                   (pc == 9'd251) ?  {5'd12,  4'd1} :
                   (pc == 9'd252) ?  {5'd0,  4'd1} :
                   (pc == 9'd253) ?  {5'd11,  4'd1} :
                   (pc == 9'd254) ?  {5'd10,  4'd1} :
                   (pc == 9'd255) ?  {5'd0,  4'd1} ://40�@�E�E�E���E�V�E�V���E
                   (pc == 9'd256) ?  {5'd8,  4'd2} :
                   (pc == 9'd257) ?  {5'd17,  4'd2} :
                   (pc == 9'd258) ?  {5'd20,  4'd1} :
                   (pc == 9'd259) ?  {5'd23,  4'd1} :
                   (pc == 9'd260) ?  {5'd0,  4'd1} :
                   (pc == 9'd261) ?  {5'd18,  4'd1} :
                   (pc == 9'd262) ?  {5'd20,  4'd1} ://41�@�\�~�\���E�t�@�\
                   (pc == 9'd263) ?  {5'd0,  4'd1} :
                   (pc == 9'd264) ?  {5'd17,  4'd1} :
                   (pc == 9'd265) ?  {5'd0,  4'd1} :
                   (pc == 9'd266) ?  {5'd13,  4'd1} :
                   (pc == 9'd267) ?  {5'd15,  4'd1} :
                   (pc == 9'd268) ?  {5'd12,  4'd1} :
                   (pc == 9'd269) ?  {5'd0,  4'd3} : //42�@�E�~�E�h���V�E�E�E (�Q�T�ڏI��)
                   (pc == 9'd270) ?  {5'd17,  4'd1} :
                   (pc == 9'd271) ?  {5'd13,  4'd1} :
                   (pc == 9'd272) ?  {5'd0,  4'd1} :
                   (pc == 9'd273) ?  {5'd8,  4'd1} :
                   (pc == 9'd274) ?  {5'd0,  4'd3} :
                   (pc == 9'd275) ?  {5'd9,  4'd1} :
                   (pc == 9'd276) ?  {5'd0,  4'd1} ://43�@�~�h�E�\�E�\
                   (pc == 9'd277) ?  {5'd10,  4'd1} :
                   (pc == 9'd278) ?  {5'd18,  4'd1} :
                   (pc == 9'd279) ?  {5'd0,  4'd1} :
                   (pc == 9'd280) ?  {5'd18,  4'd1} :
                   (pc == 9'd281) ?  {5'd10,  4'd1} :
                   (pc == 9'd282) ?  {5'd0,  4'd5} ://44�@���t�@�E�t�@��
                   (pc == 9'd283) ?  {5'd12,  4'd2} :
                   (pc == 9'd284) ?  {5'd23,  4'd2} :
                   (pc == 9'd285) ?  {5'd23,  4'd1} :
                   (pc == 9'd286) ?  {5'd23,  4'd2} :
                   (pc == 9'd287) ?  {5'd20,  4'd2} :
                   (pc == 9'd288) ?  {5'd18,  4'd1} ://45�@�V�������\�t�@
                   (pc == 9'd289) ?  {5'd17,  4'd1} :
                   (pc == 9'd290) ?  {5'd13,  4'd1} :
                   (pc == 9'd291) ?  {5'd0,  4'd1} :
                   (pc == 9'd292) ?  {5'd10,  4'd1} :
                   (pc == 9'd293) ?  {5'd8,  4'd1} :
                   (pc == 9'd294) ?  {5'd0,  4'd5} ://46�@�~�h���\
                   (pc == 9'd295) ?  {5'd17,  4'd1} :
                   (pc == 9'd296) ?  {5'd13,  4'd1} :
                   (pc == 9'd297) ?  {5'd0,  4'd1} :
                   (pc == 9'd298) ?  {5'd8,  4'd1} :
                   (pc == 9'd299) ?  {5'd0,  4'd3} :
                   (pc == 9'd300) ?  {5'd9,  4'd1} :
                   (pc == 9'd301) ?  {5'd0,  4'd1} ://47�@�~�h�E�\�E�\
                   (pc == 9'd302) ?  {5'd10,  4'd1} :
                   (pc == 9'd303) ?  {5'd18,  4'd1} :
                   (pc == 9'd304) ?  {5'd0,  4'd1} :
                   (pc == 9'd305) ?  {5'd18,  4'd1} :
                   (pc == 9'd306) ?  {5'd10,  4'd1} :
                   (pc == 9'd307) ?  {5'd0,  4'd5} ://48�@���t�@�E�t�@��
                   (pc == 9'd308) ?  {5'd12,  4'd1} :
                   (pc == 9'd309) ?  {5'd18,  4'd1} :
                   (pc == 9'd310) ?  {5'd0,  4'd1} :
                   (pc == 9'd311) ?  {5'd18,  4'd1} :
                   (pc == 9'd312) ?  {5'd18,  4'd2} :
                   (pc == 9'd313) ?  {5'd17,  4'd2} :
                   (pc == 9'd314) ?  {5'd15,  4'd1} ://49�@�V�t�@�t�@�t�@�~���h
                   (pc == 9'd315) ?  {5'd13,  4'd1} :
                   (pc == 9'd316) ?  {5'd0,  4'd13} ://50�@�h�E�E�E
                   (pc == 9'd317) ?  {5'd17,  4'd1} :
                   (pc == 9'd318) ?  {5'd13,  4'd1} :
                   (pc == 9'd319) ?  {5'd0,  4'd1} :
                   (pc == 9'd320) ?  {5'd8,  4'd1} :
                   (pc == 9'd321) ?  {5'd0,  4'd3} :
                   (pc == 9'd322) ?  {5'd9,  4'd1} :
                   (pc == 9'd323) ?  {5'd0,  4'd1} ://51�@�~�h�E�\�E�\
                   (pc == 9'd324) ?  {5'd10,  4'd1} :
                   (pc == 9'd325) ?  {5'd18,  4'd1} :
                   (pc == 9'd326) ?  {5'd0,  4'd1} :
                   (pc == 9'd327) ?  {5'd18,  4'd1} :
                   (pc == 9'd328) ?  {5'd10,  4'd1} :
                   (pc == 9'd329) ?  {5'd0,  4'd5} ://52�@���t�@�E�t�@��
                   (pc == 9'd330) ?  {5'd12,  4'd2} :
                   (pc == 9'd331) ?  {5'd23,  4'd2} :
                   (pc == 9'd332) ?  {5'd23,  4'd1} :
                   (pc == 9'd333) ?  {5'd23,  4'd2} :
                   (pc == 9'd334) ?  {5'd20,  4'd2} :
                   (pc == 9'd335) ?  {5'd18,  4'd1} ://53�@�V�������\�t�@
                   (pc == 9'd336) ?  {5'd17,  4'd1} :
                   (pc == 9'd337) ?  {5'd13,  4'd1} :
                   (pc == 9'd338) ?  {5'd0,  4'd1} :
                   (pc == 9'd339) ?  {5'd10,  4'd1} :
                   (pc == 9'd340) ?  {5'd8,  4'd1} :
                   (pc == 9'd341) ?  {5'd0,  4'd5} ://54�@�~�h���\
                   (pc == 9'd342) ?  {5'd17,  4'd1} :
                   (pc == 9'd343) ?  {5'd13,  4'd1} :
                   (pc == 9'd344) ?  {5'd0,  4'd1} :
                   (pc == 9'd345) ?  {5'd8,  4'd1} :
                   (pc == 9'd346) ?  {5'd0,  4'd3} :
                   (pc == 9'd347) ?  {5'd9,  4'd1} :
                   (pc == 9'd348) ?  {5'd0,  4'd1} ://55�@�~�h�E�\�E�\
                   (pc == 9'd349) ?  {5'd10,  4'd1} :
                   (pc == 9'd350) ?  {5'd18,  4'd1} :
                   (pc == 9'd351) ?  {5'd0,  4'd1} :
                   (pc == 9'd352) ?  {5'd18,  4'd1} :
                   (pc == 9'd353) ?  {5'd10,  4'd1} :
                   (pc == 9'd354) ?  {5'd0,  4'd5} ://56�@���t�@�E�t�@��
                   (pc == 9'd355) ?  {5'd12,  4'd1} :
                   (pc == 9'd356) ?  {5'd18,  4'd1} :
                   (pc == 9'd357) ?  {5'd0,  4'd1} :
                   (pc == 9'd358) ?  {5'd18,  4'd1} :
                   (pc == 9'd359) ?  {5'd18,  4'd2} :
                   (pc == 9'd360) ?  {5'd17,  4'd2} :
                   (pc == 9'd361) ?  {5'd15,  4'd1} ://57�@�V�t�@�t�@�t�@�~���h
                   (pc == 9'd362) ?  {5'd13,  4'd1} :
                   (pc == 9'd363) ?  {5'd0,  4'd13} ://58�@�h�E�E�E
                   (pc == 9'd364) ?  {5'd13,  4'd1} :
                   (pc == 9'd365) ?  {5'd13,  4'd1} :
                   (pc == 9'd366) ?  {5'd0,  4'd1} :
                   (pc == 9'd367) ?  {5'd13,  4'd1} :
                   (pc == 9'd368) ?  {5'd0,  4'd1} :
                   (pc == 9'd369) ?  {5'd13,  4'd1} :
                   (pc == 9'd370) ?  {5'd15,  4'd1} :
                   (pc == 9'd371) ?  {5'd0,  4'd1} ://59�@�h�h�E�h�E�h��
                   (pc == 9'd372) ?  {5'd17,  4'd1} :
                   (pc == 9'd373) ?  {5'd13,  4'd1} :
                   (pc == 9'd374) ?  {5'd0,  4'd1} :
                   (pc == 9'd375) ?  {5'd10,  4'd1} :
                   (pc == 9'd376) ?  {5'd8,  4'd1} :
                   (pc == 9'd377) ?  {5'd0,  4'd5} ://60�@�~�h���\
                   (pc == 9'd378) ?  {5'd13,  4'd1} :
                   (pc == 9'd379) ?  {5'd13,  4'd1} :
                   (pc == 9'd380) ?  {5'd0,  4'd1} :
                   (pc == 9'd381) ?  {5'd13,  4'd1} :
                   (pc == 9'd382) ?  {5'd0,  4'd1} :
                   (pc == 9'd383) ?  {5'd13,  4'd1} :
                   (pc == 9'd384) ?  {5'd15,  4'd1} :
                   (pc == 9'd385) ?  {5'd17,  4'd1} ://61�@�h�h�E�h�E�h���~
                   (pc == 9'd386) ?  {5'd0,  4'd15} ://62�@�E�E�E
                   (pc == 9'd387) ?  {5'd13,  4'd1} :
                   (pc == 9'd388) ?  {5'd13,  4'd1} :
                   (pc == 9'd389) ?  {5'd0,  4'd1} :
                   (pc == 9'd390) ?  {5'd13,  4'd1} :
                   (pc == 9'd391) ?  {5'd0,  4'd1} :
                   (pc == 9'd392) ?  {5'd13,  4'd1} :
                   (pc == 9'd393) ?  {5'd15,  4'd1} :
                   (pc == 9'd394) ?  {5'd0,  4'd1} ://63�@�h�h�E�h�E�h��
                   (pc == 9'd395) ?  {5'd17,  4'd1} :
                   (pc == 9'd396) ?  {5'd13,  4'd1} :
                   (pc == 9'd397) ?  {5'd0,  4'd1} :
                   (pc == 9'd398) ?  {5'd10,  4'd1} :
                   (pc == 9'd399) ?  {5'd8,  4'd1} :
                   (pc == 9'd400) ?  {5'd0,  4'd5} ://64�@�~�h���\
                   (pc == 9'd401)  ?  {5'd17, 4'd1} :
                   (pc == 9'd402)  ?  {5'd17, 4'd1} :
                   (pc == 9'd403)  ?  {5'd0,  4'd1} :
                   (pc == 9'd404)  ?  {5'd17, 4'd1} :
                   (pc == 9'd405)  ?  {5'd0 , 4'd1} :
                   (pc == 9'd406)  ?  {5'd13, 4'd1} :
                   (pc == 9'd407)  ?  {5'd17, 4'd1} :
                   (pc == 9'd408)  ?  {5'd0,  4'd1} ://65�@�~�~�E�~�E�h�~�E
                   (pc == 9'd409)  ?  {5'd20, 4'd1} :
                   (pc == 9'd410) ?  {5'd0,  4'd5} :
                   (pc == 9'd411) ?  {5'd8,  4'd1} :
                   (pc == 9'd412) ?  {5'd0,  4'd5} ://66�@�\�E�E�E�\�E�E�E
                   (pc == 9'd413) ?  {5'd17,  4'd1} :
                   (pc == 9'd414) ?  {5'd13,  4'd1} :
                   (pc == 9'd415) ?  {5'd0,  4'd1} :
                   (pc == 9'd416) ?  {5'd8,  4'd1} :
                   (pc == 9'd417) ?  {5'd0,  4'd3} :
                   (pc == 9'd418) ?  {5'd9,  4'd1} :
                   (pc == 9'd419) ?  {5'd0,  4'd1} ://67�@�~�h�E�\�E�\
                   (pc == 9'd420) ?  {5'd10,  4'd1} :
                   (pc == 9'd421) ?  {5'd18,  4'd1} :
                   (pc == 9'd422) ?  {5'd0,  4'd1} :
                   (pc == 9'd423) ?  {5'd18,  4'd1} :
                   (pc == 9'd424) ?  {5'd10,  4'd1} :
                   (pc == 9'd425) ?  {5'd0,  4'd5} ://68�@���t�@�E�t�@��
                   (pc == 9'd426) ?  {5'd12,  4'd2} :
                   (pc == 9'd427) ?  {5'd23,  4'd2} :
                   (pc == 9'd428) ?  {5'd23,  4'd1} :
                   (pc == 9'd429) ?  {5'd23,  4'd2} :
                   (pc == 9'd430) ?  {5'd20,  4'd2} :
                   (pc == 9'd431) ?  {5'd18,  4'd1} ://69�@�V�������\�t�@
                   (pc == 9'd432) ?  {5'd17,  4'd1} :
                   (pc == 9'd433) ?  {5'd13,  4'd1} :
                   (pc == 9'd434) ?  {5'd0,  4'd1} :
                   (pc == 9'd435) ?  {5'd10,  4'd1} :
                   (pc == 9'd436) ?  {5'd8,  4'd1} :
                   (pc == 9'd437) ?  {5'd0,  4'd5} ://70�@�~�h���\
                   (pc == 9'd438) ?  {5'd17,  4'd1} :
                   (pc == 9'd439) ?  {5'd13,  4'd1} :
                   (pc == 9'd440) ?  {5'd0,  4'd1} :
                   (pc == 9'd441) ?  {5'd8,  4'd1} :
                   (pc == 9'd442) ?  {5'd0,  4'd3} :
                   (pc == 9'd443) ?  {5'd9,  4'd1} :
                   (pc == 9'd444) ?  {5'd0,  4'd1} ://71�@�~�h�E�\�E�\
                   (pc == 9'd445) ?  {5'd10,  4'd1} :
                   (pc == 9'd446) ?  {5'd18,  4'd1} :
                   (pc == 9'd447) ?  {5'd0,  4'd1} :
                   (pc == 9'd448) ?  {5'd18,  4'd1} :
                   (pc == 9'd449) ?  {5'd10,  4'd1} :
                   (pc == 9'd450) ?  {5'd0,  4'd5} ://72�@���t�@�E�t�@��
                   (pc == 9'd451) ?  {5'd12,  4'd1} :
                   (pc == 9'd452) ?  {5'd18,  4'd1} :
                   (pc == 9'd453) ?  {5'd0,  4'd1} :
                   (pc == 9'd454) ?  {5'd18,  4'd1} :
                   (pc == 9'd455) ?  {5'd18,  4'd2} :
                   (pc == 9'd456) ?  {5'd17,  4'd2} :
                   (pc == 9'd457) ?  {5'd15,  4'd1} ://73�@�V�t�@�t�@�t�@�~���h
                   (pc == 9'd458) ?  {5'd13,  4'd1} :
                   (pc == 9'd459) ?  {5'd0,  4'd13} ://74�@�h�E�E�E
                   {5'd0, 4'd0};

    
endmodule